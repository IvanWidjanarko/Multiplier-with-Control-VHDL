LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY Multiplier_with_Control IS
	PORT
	(
		CLOCK				:	IN		BIT;
		ST					:	IN		BIT;
		MULTIPLIER		:	IN		BIT_VECTOR	(15 DOWNTO 0);
		MULTIPLICAND	:	IN		BIT_VECTOR	(15 DOWNTO 0);
		PRODUCT			:	OUT	BIT_VECTOR	(31 DOWNTO 0);
		DONE				:	INOUT	BIT
	);
END Multiplier_with_Control;

ARCHITECTURE Mul_w_Cont OF Multiplier_with_Control IS
	SIGNAL	STATE					:	INTEGER RANGE 0 TO 5;
	SIGNAL	NEXT_STATE			:	INTEGER RANGE 0 TO 5;
	SIGNAL	ACC_MULTIPLICAND	:	BIT_VECTOR	(15 DOWNTO 0);
	SIGNAL	ACC_MULTIPLIER		:	BIT_VECTOR	(15 DOWNTO 0);
	SIGNAL	ADSH					:	BIT;
	SIGNAL	SH						:	BIT;
	SIGNAL	LOAD					:	BIT;
	SIGNAL	CM						:	BIT;
	ALIAS		M						:	BIT	IS	ACC_MULTIPLIER(0);
	
	FUNCTION ADD4 (REG1,REG2: BIT_VECTOR(15 DOWNTO 0);CARRY: BIT) 
	RETURN BIT_VECTOR IS
		VARIABLE COUT: BIT:='0';
		VARIABLE CIN: BIT:=CARRY;
		VARIABLE RETVAL: BIT_VECTOR(16 DOWNTO 0):="00000000000000000";
		BEGIN
		LP1: FOR I IN 0 TO 3 LOOP
			COUT :=(REG1(I) AND REG2(I)) OR ( REG1(I) AND CIN) OR 
						(REG2(I) AND CIN );
			RETVAL(I) := REG1(I) XOR REG2(I) XOR CIN;
			CIN := COUT; 
		END LOOP LP1;
		RETVAL(4):=COUT;
		RETURN RETVAL;
	END ADD4;

BEGIN

	Multiplier_2s_Complement : PROCESS
	
	VARIABLE	ADDOUT				:	BIT_VECTOR	(16 DOWNTO 0);
	
	BEGIN
	
		LOAD	<=	'0';
		ADSH	<=	'0';
		SH		<=	'0';
		CM		<=	'0';
		DONE	<=	'0';
		
		CASE	STATE	IS
			WHEN	0	=>
				IF ST='1' THEN
					LOAD			<=	'1';
					NEXT_STATE	<=	1;
				END IF;
			WHEN 1 | 2 | 3	=>
				IF M = '1' THEN
					ADSH		<=	'1';
				ELSE
					SH			<= '1';
				END IF;
				NEXT_STATE	<=	STATE + 1;
			WHEN 4	=>
				IF M = '1'THEN
					CM		<=	'1';
					ADSH	<=	'1';
				ELSE
					SH		<=	'1';
				END IF;
				NEXT_STATE	<= 5;
			WHEN 5	=>
				DONE			<=	'1';
				NEXT_sTATE	<=	0;
		END CASE;
	
		WAIT UNTIL CLOCK ='1';
		
		IF CM = '0' THEN
			ADDOUT	:=	ADD4(ACC_MULTIPLICAND,MULTIPLICAND,'0');
		ELSE
			ADDOUT	:=	ADD4(ACC_MULTIPLICAND, NOT MULTIPLICAND,'1');
		END IF;
		
		IF LOAD = '1'THEN
			ACC_MULTIPLICAND	<=	"0000000000000000";
			ACC_MULTIPLIER		<=	MULTIPLIER;
		END IF;
		
		IF ADSH = '1'THEN
			ACC_MULTIPLICAND	<=	(MULTIPLICAND(15) XOR CM) & ADDOUT(15 DOWNTO 1);
			ACC_MULTIPLIER		<= ADDOUT(0) & ACC_MULTIPLIER(15 DOWNTO 1);
		END IF;
		
		IF SH = '1'THEN
			ACC_MULTIPLICAND	<= ACC_MULTIPLICAND(15) & ACC_MULTIPLICAND(15 DOWNTO 1);
			ACC_MULTIPLICAND	<=	ACC_MULTIPLICAND(0) & ACC_MULTIPLIER(15 DOWNTO 1);
		END IF;
		
		IF DONE = '1' THEN
			Product <= ACC_MULTIPLICAND(15 downto 0) & ACC_MULTIPLIER;
		END IF;
		
		STATE	<=	NEXT_STATE;
	
	END PROCESS Multiplier_2s_Complement;
	
END Mul_w_Cont;